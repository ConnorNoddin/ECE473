// Connor Noddin
// ECE 473
// ID_EX Block
// 10/07/2023

module EX_MEM(
	input wire clock,
	input wire reset,
	input wire [31:0] D1_IN,
	input wire [31:0] D2_IN,
	input wire [4:0] RD_IN,
	output reg [31:0] D1_MEM,
	output reg [31:0] D2_MEM,
	output reg [4:0] RD_MEM);
	
	// Write data on positive edge or reset
	always @(posedge clock or posedge reset) begin
		if(reset == 1'b1) begin
			D1_MEM <= 32'd0;
			D2_MEM <= 32'd0;
			RD_MEM <= 5'd0;
		end else begin
			D1_MEM <= D1_IN;
			D2_MEM <= D2_IN;
			RD_MEM <= RD_IN;
		end
	end
	
endmodule

